-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Array_pkg.all;
use work.mmio_pkg.all;

entity Kernel_Nucleus is
  generic (
    INDEX_WIDTH                       : integer := 32;
    TAG_WIDTH                         : integer := 1;
    STRINGWRITE_STRING_BUS_ADDR_WIDTH : integer := 64
  );
  port (
    kcd_clk                         : in  std_logic;
    kcd_reset                       : in  std_logic;
    mmio_awvalid                    : in  std_logic;
    mmio_awready                    : out std_logic;
    mmio_awaddr                     : in  std_logic_vector(31 downto 0);
    mmio_wvalid                     : in  std_logic;
    mmio_wready                     : out std_logic;
    mmio_wdata                      : in  std_logic_vector(31 downto 0);
    mmio_wstrb                      : in  std_logic_vector(3 downto 0);
    mmio_bvalid                     : out std_logic;
    mmio_bready                     : in  std_logic;
    mmio_bresp                      : out std_logic_vector(1 downto 0);
    mmio_arvalid                    : in  std_logic;
    mmio_arready                    : out std_logic;
    mmio_araddr                     : in  std_logic_vector(31 downto 0);
    mmio_rvalid                     : out std_logic;
    mmio_rready                     : in  std_logic;
    mmio_rdata                      : out std_logic_vector(31 downto 0);
    mmio_rresp                      : out std_logic_vector(1 downto 0);
    StringWrite_String_valid        : out std_logic;
    StringWrite_String_ready        : in  std_logic;
    StringWrite_String_dvalid       : out std_logic;
    StringWrite_String_last         : out std_logic;
    StringWrite_String_length       : out std_logic_vector(31 downto 0);
    StringWrite_String_count        : out std_logic_vector(0 downto 0);
    StringWrite_String_chars_valid  : out std_logic;
    StringWrite_String_chars_ready  : in  std_logic;
    StringWrite_String_chars_dvalid : out std_logic;
    StringWrite_String_chars_last   : out std_logic;
    StringWrite_String_chars        : out std_logic_vector(511 downto 0);
    StringWrite_String_chars_count  : out std_logic_vector(6 downto 0);
    StringWrite_String_unl_valid    : in  std_logic;
    StringWrite_String_unl_ready    : out std_logic;
    StringWrite_String_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    StringWrite_String_cmd_valid    : out std_logic;
    StringWrite_String_cmd_ready    : in  std_logic;
    StringWrite_String_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    StringWrite_String_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    StringWrite_String_cmd_ctrl     : out std_logic_vector(STRINGWRITE_STRING_BUS_ADDR_WIDTH*2-1 downto 0);
    StringWrite_String_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0)
  );
end entity;

architecture Implementation of Kernel_Nucleus is
  component Kernel is
    generic (
      INDEX_WIDTH : integer := 32;
      TAG_WIDTH   : integer := 1
    );
    port (
      kcd_clk                         : in  std_logic;
      kcd_reset                       : in  std_logic;
      StringWrite_String_valid        : out std_logic;
      StringWrite_String_ready        : in  std_logic;
      StringWrite_String_dvalid       : out std_logic;
      StringWrite_String_last         : out std_logic;
      StringWrite_String_length       : out std_logic_vector(31 downto 0);
      StringWrite_String_count        : out std_logic_vector(0 downto 0);
      StringWrite_String_chars_valid  : out std_logic;
      StringWrite_String_chars_ready  : in  std_logic;
      StringWrite_String_chars_dvalid : out std_logic;
      StringWrite_String_chars_last   : out std_logic;
      StringWrite_String_chars        : out std_logic_vector(511 downto 0);
      StringWrite_String_chars_count  : out std_logic_vector(6 downto 0);
      StringWrite_String_unl_valid    : in  std_logic;
      StringWrite_String_unl_ready    : out std_logic;
      StringWrite_String_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      StringWrite_String_cmd_valid    : out std_logic;
      StringWrite_String_cmd_ready    : in  std_logic;
      StringWrite_String_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      StringWrite_String_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      StringWrite_String_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      start                           : in  std_logic;
      stop                            : in  std_logic;
      reset                           : in  std_logic;
      idle                            : out std_logic;
      busy                            : out std_logic;
      done                            : out std_logic;
      result                          : out std_logic_vector(63 downto 0);
      StringWrite_firstidx            : in  std_logic_vector(31 downto 0);
      StringWrite_lastidx             : in  std_logic_vector(31 downto 0);
      strlen_min                      : in  std_logic_vector(31 downto 0);
      strlen_mask                     : in  std_logic_vector(31 downto 0)
    );
  end component;

  signal Kernel_inst_kcd_clk                                   : std_logic;
  signal Kernel_inst_kcd_reset                                 : std_logic;

  signal Kernel_inst_StringWrite_String_valid                  : std_logic;
  signal Kernel_inst_StringWrite_String_ready                  : std_logic;
  signal Kernel_inst_StringWrite_String_dvalid                 : std_logic;
  signal Kernel_inst_StringWrite_String_last                   : std_logic;
  signal Kernel_inst_StringWrite_String_length                 : std_logic_vector(31 downto 0);
  signal Kernel_inst_StringWrite_String_count                  : std_logic_vector(0 downto 0);
  signal Kernel_inst_StringWrite_String_chars_valid            : std_logic;
  signal Kernel_inst_StringWrite_String_chars_ready            : std_logic;
  signal Kernel_inst_StringWrite_String_chars_dvalid           : std_logic;
  signal Kernel_inst_StringWrite_String_chars_last             : std_logic;
  signal Kernel_inst_StringWrite_String_chars                  : std_logic_vector(511 downto 0);
  signal Kernel_inst_StringWrite_String_chars_count            : std_logic_vector(6 downto 0);

  signal Kernel_inst_StringWrite_String_unl_valid              : std_logic;
  signal Kernel_inst_StringWrite_String_unl_ready              : std_logic;
  signal Kernel_inst_StringWrite_String_unl_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_StringWrite_String_cmd_valid              : std_logic;
  signal Kernel_inst_StringWrite_String_cmd_ready              : std_logic;
  signal Kernel_inst_StringWrite_String_cmd_firstIdx           : std_logic_vector(31 downto 0);
  signal Kernel_inst_StringWrite_String_cmd_lastIdx            : std_logic_vector(31 downto 0);
  signal Kernel_inst_StringWrite_String_cmd_tag                : std_logic_vector(0 downto 0);

  signal Kernel_inst_start                                     : std_logic;
  signal Kernel_inst_stop                                      : std_logic;
  signal Kernel_inst_reset                                     : std_logic;
  signal Kernel_inst_idle                                      : std_logic;
  signal Kernel_inst_busy                                      : std_logic;
  signal Kernel_inst_done                                      : std_logic;
  signal Kernel_inst_result                                    : std_logic_vector(63 downto 0);
  signal Kernel_inst_StringWrite_firstidx                      : std_logic_vector(31 downto 0);
  signal Kernel_inst_StringWrite_lastidx                       : std_logic_vector(31 downto 0);
  signal Kernel_inst_strlen_min                                : std_logic_vector(31 downto 0);
  signal Kernel_inst_strlen_mask                               : std_logic_vector(31 downto 0);
  signal mmio_inst_kcd_clk                                     : std_logic;
  signal mmio_inst_kcd_reset                                   : std_logic;

  signal mmio_inst_f_start_data                                : std_logic;
  signal mmio_inst_f_stop_data                                 : std_logic;
  signal mmio_inst_f_reset_data                                : std_logic;
  signal mmio_inst_f_idle_write_data                           : std_logic;
  signal mmio_inst_f_busy_write_data                           : std_logic;
  signal mmio_inst_f_done_write_data                           : std_logic;
  signal mmio_inst_f_result_write_data                         : std_logic_vector(63 downto 0);
  signal mmio_inst_f_StringWrite_firstidx_data                 : std_logic_vector(31 downto 0);
  signal mmio_inst_f_StringWrite_lastidx_data                  : std_logic_vector(31 downto 0);
  signal mmio_inst_f_StringWrite_String_offsets_data           : std_logic_vector(63 downto 0);
  signal mmio_inst_f_StringWrite_String_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_strlen_min_data                           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_strlen_mask_data                          : std_logic_vector(31 downto 0);
  signal mmio_inst_f_Profile_enable_data                       : std_logic;
  signal mmio_inst_f_Profile_clear_data                        : std_logic;
  signal mmio_inst_mmio_awvalid                                : std_logic;
  signal mmio_inst_mmio_awready                                : std_logic;
  signal mmio_inst_mmio_awaddr                                 : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_wvalid                                 : std_logic;
  signal mmio_inst_mmio_wready                                 : std_logic;
  signal mmio_inst_mmio_wdata                                  : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_wstrb                                  : std_logic_vector(3 downto 0);
  signal mmio_inst_mmio_bvalid                                 : std_logic;
  signal mmio_inst_mmio_bready                                 : std_logic;
  signal mmio_inst_mmio_bresp                                  : std_logic_vector(1 downto 0);
  signal mmio_inst_mmio_arvalid                                : std_logic;
  signal mmio_inst_mmio_arready                                : std_logic;
  signal mmio_inst_mmio_araddr                                 : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_rvalid                                 : std_logic;
  signal mmio_inst_mmio_rready                                 : std_logic;
  signal mmio_inst_mmio_rdata                                  : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_rresp                                  : std_logic_vector(1 downto 0);

  signal StringWrite_String_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal StringWrite_String_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal StringWrite_String_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal StringWrite_String_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal StringWrite_String_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal StringWrite_String_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal StringWrite_String_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal StringWrite_String_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal StringWrite_String_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal StringWrite_String_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(2*STRINGWRITE_STRING_BUS_ADDR_WIDTH-1 downto 0);
  signal StringWrite_String_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal StringWrite_String_cmd_accm_inst_ctrl : std_logic_vector(2*STRINGWRITE_STRING_BUS_ADDR_WIDTH-1 downto 0);

begin
  Kernel_inst : Kernel
    generic map (
      INDEX_WIDTH => 32,
      TAG_WIDTH   => 1
    )
    port map (
      kcd_clk                         => Kernel_inst_kcd_clk,
      kcd_reset                       => Kernel_inst_kcd_reset,
      StringWrite_String_valid        => Kernel_inst_StringWrite_String_valid,
      StringWrite_String_ready        => Kernel_inst_StringWrite_String_ready,
      StringWrite_String_dvalid       => Kernel_inst_StringWrite_String_dvalid,
      StringWrite_String_last         => Kernel_inst_StringWrite_String_last,
      StringWrite_String_length       => Kernel_inst_StringWrite_String_length,
      StringWrite_String_count        => Kernel_inst_StringWrite_String_count,
      StringWrite_String_chars_valid  => Kernel_inst_StringWrite_String_chars_valid,
      StringWrite_String_chars_ready  => Kernel_inst_StringWrite_String_chars_ready,
      StringWrite_String_chars_dvalid => Kernel_inst_StringWrite_String_chars_dvalid,
      StringWrite_String_chars_last   => Kernel_inst_StringWrite_String_chars_last,
      StringWrite_String_chars        => Kernel_inst_StringWrite_String_chars,
      StringWrite_String_chars_count  => Kernel_inst_StringWrite_String_chars_count,
      StringWrite_String_unl_valid    => Kernel_inst_StringWrite_String_unl_valid,
      StringWrite_String_unl_ready    => Kernel_inst_StringWrite_String_unl_ready,
      StringWrite_String_unl_tag      => Kernel_inst_StringWrite_String_unl_tag,
      StringWrite_String_cmd_valid    => Kernel_inst_StringWrite_String_cmd_valid,
      StringWrite_String_cmd_ready    => Kernel_inst_StringWrite_String_cmd_ready,
      StringWrite_String_cmd_firstIdx => Kernel_inst_StringWrite_String_cmd_firstIdx,
      StringWrite_String_cmd_lastIdx  => Kernel_inst_StringWrite_String_cmd_lastIdx,
      StringWrite_String_cmd_tag      => Kernel_inst_StringWrite_String_cmd_tag,
      start                           => Kernel_inst_start,
      stop                            => Kernel_inst_stop,
      reset                           => Kernel_inst_reset,
      idle                            => Kernel_inst_idle,
      busy                            => Kernel_inst_busy,
      done                            => Kernel_inst_done,
      result                          => Kernel_inst_result,
      StringWrite_firstidx            => Kernel_inst_StringWrite_firstidx,
      StringWrite_lastidx             => Kernel_inst_StringWrite_lastidx,
      strlen_min                      => Kernel_inst_strlen_min,
      strlen_mask                     => Kernel_inst_strlen_mask
    );

  mmio_inst : mmio
    port map (
      kcd_clk                           => mmio_inst_kcd_clk,
      kcd_reset                         => mmio_inst_kcd_reset,
      f_start_data                      => mmio_inst_f_start_data,
      f_stop_data                       => mmio_inst_f_stop_data,
      f_reset_data                      => mmio_inst_f_reset_data,
      f_idle_write_data                 => mmio_inst_f_idle_write_data,
      f_busy_write_data                 => mmio_inst_f_busy_write_data,
      f_done_write_data                 => mmio_inst_f_done_write_data,
      f_result_write_data               => mmio_inst_f_result_write_data,
      f_StringWrite_firstidx_data       => mmio_inst_f_StringWrite_firstidx_data,
      f_StringWrite_lastidx_data        => mmio_inst_f_StringWrite_lastidx_data,
      f_StringWrite_String_offsets_data => mmio_inst_f_StringWrite_String_offsets_data,
      f_StringWrite_String_values_data  => mmio_inst_f_StringWrite_String_values_data,
      f_strlen_min_data                 => mmio_inst_f_strlen_min_data,
      f_strlen_mask_data                => mmio_inst_f_strlen_mask_data,
      mmio_awvalid                      => mmio_inst_mmio_awvalid,
      mmio_awready                      => mmio_inst_mmio_awready,
      mmio_awaddr                       => mmio_inst_mmio_awaddr,
      mmio_wvalid                       => mmio_inst_mmio_wvalid,
      mmio_wready                       => mmio_inst_mmio_wready,
      mmio_wdata                        => mmio_inst_mmio_wdata,
      mmio_wstrb                        => mmio_inst_mmio_wstrb,
      mmio_bvalid                       => mmio_inst_mmio_bvalid,
      mmio_bready                       => mmio_inst_mmio_bready,
      mmio_bresp                        => mmio_inst_mmio_bresp,
      mmio_arvalid                      => mmio_inst_mmio_arvalid,
      mmio_arready                      => mmio_inst_mmio_arready,
      mmio_araddr                       => mmio_inst_mmio_araddr,
      mmio_rvalid                       => mmio_inst_mmio_rvalid,
      mmio_rready                       => mmio_inst_mmio_rready,
      mmio_rdata                        => mmio_inst_mmio_rdata,
      mmio_rresp                        => mmio_inst_mmio_rresp
    );

  StringWrite_String_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => STRINGWRITE_STRING_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => StringWrite_String_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => StringWrite_String_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => StringWrite_String_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => StringWrite_String_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => StringWrite_String_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => StringWrite_String_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => StringWrite_String_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => StringWrite_String_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => StringWrite_String_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => StringWrite_String_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => StringWrite_String_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => StringWrite_String_cmd_accm_inst_ctrl
    );

  StringWrite_String_valid                           <= Kernel_inst_StringWrite_String_valid;
  Kernel_inst_StringWrite_String_ready               <= StringWrite_String_ready;
  StringWrite_String_dvalid                          <= Kernel_inst_StringWrite_String_dvalid;
  StringWrite_String_last                            <= Kernel_inst_StringWrite_String_last;
  StringWrite_String_length                          <= Kernel_inst_StringWrite_String_length;
  StringWrite_String_count                           <= Kernel_inst_StringWrite_String_count;
  StringWrite_String_chars_valid                     <= Kernel_inst_StringWrite_String_chars_valid;
  Kernel_inst_StringWrite_String_chars_ready         <= StringWrite_String_chars_ready;
  StringWrite_String_chars_dvalid                    <= Kernel_inst_StringWrite_String_chars_dvalid;
  StringWrite_String_chars_last                      <= Kernel_inst_StringWrite_String_chars_last;
  StringWrite_String_chars                           <= Kernel_inst_StringWrite_String_chars;
  StringWrite_String_chars_count                     <= Kernel_inst_StringWrite_String_chars_count;

  StringWrite_String_cmd_valid                       <= StringWrite_String_cmd_accm_inst_nucleus_cmd_valid;
  StringWrite_String_cmd_accm_inst_nucleus_cmd_ready <= StringWrite_String_cmd_ready;
  StringWrite_String_cmd_firstIdx                    <= StringWrite_String_cmd_accm_inst_nucleus_cmd_firstIdx;
  StringWrite_String_cmd_lastIdx                     <= StringWrite_String_cmd_accm_inst_nucleus_cmd_lastIdx;
  StringWrite_String_cmd_ctrl                        <= StringWrite_String_cmd_accm_inst_nucleus_cmd_ctrl;
  StringWrite_String_cmd_tag                         <= StringWrite_String_cmd_accm_inst_nucleus_cmd_tag;

  Kernel_inst_kcd_clk                                  <= kcd_clk;
  Kernel_inst_kcd_reset                                <= kcd_reset;

  Kernel_inst_StringWrite_String_unl_valid             <= StringWrite_String_unl_valid;
  StringWrite_String_unl_ready                         <= Kernel_inst_StringWrite_String_unl_ready;
  Kernel_inst_StringWrite_String_unl_tag               <= StringWrite_String_unl_tag;

  Kernel_inst_start                                    <= mmio_inst_f_start_data;
  Kernel_inst_stop                                     <= mmio_inst_f_stop_data;
  Kernel_inst_reset                                    <= mmio_inst_f_reset_data;
  Kernel_inst_StringWrite_firstidx                     <= mmio_inst_f_StringWrite_firstidx_data;
  Kernel_inst_StringWrite_lastidx                      <= mmio_inst_f_StringWrite_lastidx_data;
  Kernel_inst_strlen_min                               <= mmio_inst_f_strlen_min_data;
  Kernel_inst_strlen_mask                              <= mmio_inst_f_strlen_mask_data;
  mmio_inst_kcd_clk                                    <= kcd_clk;
  mmio_inst_kcd_reset                                  <= kcd_reset;

  mmio_inst_f_idle_write_data                          <= Kernel_inst_idle;
  mmio_inst_f_busy_write_data                          <= Kernel_inst_busy;
  mmio_inst_f_done_write_data                          <= Kernel_inst_done;
  mmio_inst_f_result_write_data                        <= Kernel_inst_result;
  mmio_inst_mmio_awvalid                               <= mmio_awvalid;
  mmio_awready                                         <= mmio_inst_mmio_awready;
  mmio_inst_mmio_awaddr                                <= mmio_awaddr;
  mmio_inst_mmio_wvalid                                <= mmio_wvalid;
  mmio_wready                                          <= mmio_inst_mmio_wready;
  mmio_inst_mmio_wdata                                 <= mmio_wdata;
  mmio_inst_mmio_wstrb                                 <= mmio_wstrb;
  mmio_bvalid                                          <= mmio_inst_mmio_bvalid;
  mmio_inst_mmio_bready                                <= mmio_bready;
  mmio_bresp                                           <= mmio_inst_mmio_bresp;
  mmio_inst_mmio_arvalid                               <= mmio_arvalid;
  mmio_arready                                         <= mmio_inst_mmio_arready;
  mmio_inst_mmio_araddr                                <= mmio_araddr;
  mmio_rvalid                                          <= mmio_inst_mmio_rvalid;
  mmio_inst_mmio_rready                                <= mmio_rready;
  mmio_rdata                                           <= mmio_inst_mmio_rdata;
  mmio_rresp                                           <= mmio_inst_mmio_rresp;

  StringWrite_String_cmd_accm_inst_kernel_cmd_valid    <= Kernel_inst_StringWrite_String_cmd_valid;
  Kernel_inst_StringWrite_String_cmd_ready             <= StringWrite_String_cmd_accm_inst_kernel_cmd_ready;
  StringWrite_String_cmd_accm_inst_kernel_cmd_firstIdx <= Kernel_inst_StringWrite_String_cmd_firstIdx;
  StringWrite_String_cmd_accm_inst_kernel_cmd_lastIdx  <= Kernel_inst_StringWrite_String_cmd_lastIdx;
  StringWrite_String_cmd_accm_inst_kernel_cmd_tag      <= Kernel_inst_StringWrite_String_cmd_tag;

  StringWrite_String_cmd_accm_inst_ctrl(63 downto 0)   <= mmio_inst_f_StringWrite_String_offsets_data;
  StringWrite_String_cmd_accm_inst_ctrl(127 downto 64) <= mmio_inst_f_StringWrite_String_values_data;

end architecture;
