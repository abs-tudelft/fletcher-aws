-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Array_pkg.all;

entity Kernel_StringWrite is
  generic (
    INDEX_WIDTH                           : integer := 32;
    TAG_WIDTH                             : integer := 1;
    STRINGWRITE_STRING_BUS_ADDR_WIDTH     : integer := 64;
    STRINGWRITE_STRING_BUS_DATA_WIDTH     : integer := 512;
    STRINGWRITE_STRING_BUS_LEN_WIDTH      : integer := 8;
    STRINGWRITE_STRING_BUS_BURST_STEP_LEN : integer := 1;
    STRINGWRITE_STRING_BUS_BURST_MAX_LEN  : integer := 16
  );
  port (
    bcd_clk                            : in  std_logic;
    bcd_reset                          : in  std_logic;
    kcd_clk                            : in  std_logic;
    kcd_reset                          : in  std_logic;
    StringWrite_String_valid           : in  std_logic;
    StringWrite_String_ready           : out std_logic;
    StringWrite_String_dvalid          : in  std_logic;
    StringWrite_String_last            : in  std_logic;
    StringWrite_String_length          : in  std_logic_vector(31 downto 0);
    StringWrite_String_count           : in  std_logic_vector(0 downto 0);
    StringWrite_String_chars_valid     : in  std_logic;
    StringWrite_String_chars_ready     : out std_logic;
    StringWrite_String_chars_dvalid    : in  std_logic;
    StringWrite_String_chars_last      : in  std_logic;
    StringWrite_String_chars           : in  std_logic_vector(511 downto 0);
    StringWrite_String_chars_count     : in  std_logic_vector(6 downto 0);
    StringWrite_String_bus_wreq_valid  : out std_logic;
    StringWrite_String_bus_wreq_ready  : in  std_logic;
    StringWrite_String_bus_wreq_addr   : out std_logic_vector(STRINGWRITE_STRING_BUS_ADDR_WIDTH-1 downto 0);
    StringWrite_String_bus_wreq_len    : out std_logic_vector(STRINGWRITE_STRING_BUS_LEN_WIDTH-1 downto 0);
    StringWrite_String_bus_wdat_valid  : out std_logic;
    StringWrite_String_bus_wdat_ready  : in  std_logic;
    StringWrite_String_bus_wdat_data   : out std_logic_vector(STRINGWRITE_STRING_BUS_DATA_WIDTH-1 downto 0);
    StringWrite_String_bus_wdat_strobe : out std_logic_vector(STRINGWRITE_STRING_BUS_DATA_WIDTH/8-1 downto 0);
    StringWrite_String_bus_wdat_last   : out std_logic;
    StringWrite_String_cmd_valid       : in  std_logic;
    StringWrite_String_cmd_ready       : out std_logic;
    StringWrite_String_cmd_firstIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    StringWrite_String_cmd_lastIdx     : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    StringWrite_String_cmd_ctrl        : in  std_logic_vector(STRINGWRITE_STRING_BUS_ADDR_WIDTH*2-1 downto 0);
    StringWrite_String_cmd_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    StringWrite_String_unl_valid       : out std_logic;
    StringWrite_String_unl_ready       : in  std_logic;
    StringWrite_String_unl_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0)
  );
end entity;

architecture Implementation of Kernel_StringWrite is
  signal String_inst_bcd_clk         : std_logic;
  signal String_inst_bcd_reset       : std_logic;

  signal String_inst_kcd_clk         : std_logic;
  signal String_inst_kcd_reset       : std_logic;

  signal String_inst_cmd_valid       : std_logic;
  signal String_inst_cmd_ready       : std_logic;
  signal String_inst_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal String_inst_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal String_inst_cmd_ctrl        : std_logic_vector(STRINGWRITE_STRING_BUS_ADDR_WIDTH*2-1 downto 0);
  signal String_inst_cmd_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal String_inst_unl_valid       : std_logic;
  signal String_inst_unl_ready       : std_logic;
  signal String_inst_unl_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal String_inst_bus_wreq_valid  : std_logic;
  signal String_inst_bus_wreq_ready  : std_logic;
  signal String_inst_bus_wreq_addr   : std_logic_vector(STRINGWRITE_STRING_BUS_ADDR_WIDTH-1 downto 0);
  signal String_inst_bus_wreq_len    : std_logic_vector(STRINGWRITE_STRING_BUS_LEN_WIDTH-1 downto 0);
  signal String_inst_bus_wdat_valid  : std_logic;
  signal String_inst_bus_wdat_ready  : std_logic;
  signal String_inst_bus_wdat_data   : std_logic_vector(STRINGWRITE_STRING_BUS_DATA_WIDTH-1 downto 0);
  signal String_inst_bus_wdat_strobe : std_logic_vector(STRINGWRITE_STRING_BUS_DATA_WIDTH/8-1 downto 0);
  signal String_inst_bus_wdat_last   : std_logic;

  signal String_inst_in_valid        : std_logic_vector(1 downto 0);
  signal String_inst_in_ready        : std_logic_vector(1 downto 0);
  signal String_inst_in_data         : std_logic_vector(551 downto 0);
  signal String_inst_in_dvalid       : std_logic_vector(1 downto 0);
  signal String_inst_in_last         : std_logic_vector(1 downto 0);

begin
  String_inst : ArrayWriter
    generic map (
      BUS_ADDR_WIDTH     => STRINGWRITE_STRING_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => STRINGWRITE_STRING_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => STRINGWRITE_STRING_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => STRINGWRITE_STRING_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => STRINGWRITE_STRING_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "listprim(8;epc=64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk         => String_inst_bcd_clk,
      bcd_reset       => String_inst_bcd_reset,
      kcd_clk         => String_inst_kcd_clk,
      kcd_reset       => String_inst_kcd_reset,
      cmd_valid       => String_inst_cmd_valid,
      cmd_ready       => String_inst_cmd_ready,
      cmd_firstIdx    => String_inst_cmd_firstIdx,
      cmd_lastIdx     => String_inst_cmd_lastIdx,
      cmd_ctrl        => String_inst_cmd_ctrl,
      cmd_tag         => String_inst_cmd_tag,
      unl_valid       => String_inst_unl_valid,
      unl_ready       => String_inst_unl_ready,
      unl_tag         => String_inst_unl_tag,
      bus_wreq_valid  => String_inst_bus_wreq_valid,
      bus_wreq_ready  => String_inst_bus_wreq_ready,
      bus_wreq_addr   => String_inst_bus_wreq_addr,
      bus_wreq_len    => String_inst_bus_wreq_len,
      bus_wdat_valid  => String_inst_bus_wdat_valid,
      bus_wdat_ready  => String_inst_bus_wdat_ready,
      bus_wdat_data   => String_inst_bus_wdat_data,
      bus_wdat_strobe => String_inst_bus_wdat_strobe,
      bus_wdat_last   => String_inst_bus_wdat_last,
      in_valid        => String_inst_in_valid,
      in_ready        => String_inst_in_ready,
      in_data         => String_inst_in_data,
      in_dvalid       => String_inst_in_dvalid,
      in_last         => String_inst_in_last
    );

  StringWrite_String_bus_wreq_valid  <= String_inst_bus_wreq_valid;
  String_inst_bus_wreq_ready         <= StringWrite_String_bus_wreq_ready;
  StringWrite_String_bus_wreq_addr   <= String_inst_bus_wreq_addr;
  StringWrite_String_bus_wreq_len    <= String_inst_bus_wreq_len;
  StringWrite_String_bus_wdat_valid  <= String_inst_bus_wdat_valid;
  String_inst_bus_wdat_ready         <= StringWrite_String_bus_wdat_ready;
  StringWrite_String_bus_wdat_data   <= String_inst_bus_wdat_data;
  StringWrite_String_bus_wdat_strobe <= String_inst_bus_wdat_strobe;
  StringWrite_String_bus_wdat_last   <= String_inst_bus_wdat_last;

  StringWrite_String_unl_valid       <= String_inst_unl_valid;
  String_inst_unl_ready              <= StringWrite_String_unl_ready;
  StringWrite_String_unl_tag         <= String_inst_unl_tag;

  String_inst_bcd_clk                 <= bcd_clk;
  String_inst_bcd_reset               <= bcd_reset;

  String_inst_kcd_clk                 <= kcd_clk;
  String_inst_kcd_reset               <= kcd_reset;

  String_inst_cmd_valid               <= StringWrite_String_cmd_valid;
  StringWrite_String_cmd_ready        <= String_inst_cmd_ready;
  String_inst_cmd_firstIdx            <= StringWrite_String_cmd_firstIdx;
  String_inst_cmd_lastIdx             <= StringWrite_String_cmd_lastIdx;
  String_inst_cmd_ctrl                <= StringWrite_String_cmd_ctrl;
  String_inst_cmd_tag                 <= StringWrite_String_cmd_tag;

  String_inst_in_valid(0)             <= StringWrite_String_valid;
  String_inst_in_valid(1)             <= StringWrite_String_chars_valid;
  StringWrite_String_ready            <= String_inst_in_ready(0);
  StringWrite_String_chars_ready      <= String_inst_in_ready(1);
  String_inst_in_data(31 downto 0)    <= StringWrite_String_length;
  String_inst_in_data(32 downto 32)   <= StringWrite_String_count;
  String_inst_in_data(544 downto 33)  <= StringWrite_String_chars;
  String_inst_in_data(551 downto 545) <= StringWrite_String_chars_count;
  String_inst_in_dvalid(0)            <= StringWrite_String_dvalid;
  String_inst_in_dvalid(1)            <= StringWrite_String_chars_dvalid;
  String_inst_in_last(0)              <= StringWrite_String_last;
  String_inst_in_last(1)              <= StringWrite_String_chars_last;

end architecture;
